** Profile: "SCHEMATIC1-12V_Boost_Converter_Sim2"  [ C:\Users\carri\OneDrive\Desktop\Master's Thesis\AtInverter\sims\12V_Boost_Converter-PSpiceFiles\SCHEMATIC1\12V_Boost_Converter_Sim2.sim ] 

** Creating circuit file "12V_Boost_Converter_Sim2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3000ns 0 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
